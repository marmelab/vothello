module othello

struct Player {
	pub mut:
		celltype CellType
}